* Design:	XOR
* Created:	"Mon Dec 9 2024"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"Calibre xACT 3D"
* Version:	"v2017.4_19.14"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

* .include "XOR.pex.netlist.pex"

* Start of included file XOR.pex.netlist.pex

.subckt PM_XOR%NET16 VSS! 6 7 3 1
c1 1 VSS! 0.00524342f $X=0.432 $Y=0.0895
c2 3 VSS! 0.00337254f $X=0.4175 $Y=0.0895
r1 7 5 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.4493 $Y=0.0895 $X2=0.4465 $Y2=0.0895
r2 1 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.432 $Y=0.0895 $X2=0.4465 $Y2=0.0895
r3 3 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.4175 $Y=0.0895 $X2=0.432 $Y2=0.0895
r4 6 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.4146 $Y=0.0895 $X2=0.4175 $Y2=0.0895
.ends

.subckt PM_XOR%B VSS! 33 16 20 44 47 11 2 1 8 7 13 6 5 12 9 10
c1 1 VSS! 0.0039654f $X=0.135 $Y=0.157
c2 2 VSS! 0.00359782f $X=0.405 $Y=0.157
c3 5 VSS! 0.0835408f $X=0.135 $Y=0.157
c4 6 VSS! 0.0802712f $X=0.405 $Y=0.0465
c5 7 VSS! 0.000792401f $X=0.135 $Y=0.1455
c6 8 VSS! 0.000528513f $X=0.405 $Y=0.1455
c7 9 VSS! 0.0027412f $X=0.135 $Y=0.058
c8 10 VSS! 0.00285365f $X=0.405 $Y=0.058
c9 11 VSS! 0.0032834f $X=0.135 $Y=0.105
c10 12 VSS! 0.0179928f $X=0.378 $Y=0.058
c11 13 VSS! 0.0047868f $X=0.405 $Y=0.1455
r1 47 46 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.135 $Y=0.2245 $X2=0.135 $Y2=0.1755
r2 44 45 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.135 $Y=0.0895 $X2=0.135 $Y2=0.1385
r3 5 45 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.135 $Y=0.157 $X2=0.135 $Y2=0.1385
r4 5 46 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.135 $Y=0.157 $X2=0.135 $Y2=0.1755
r5 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.135
+ $Y=0.157 $X2=0.135 $Y2=0.157
r6 1 5 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08 $X=0.135
+ $Y=0.157 $X2=0.135 $Y2=0.157
r7 7 39 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1455 $X2=0.135 $Y2=0.157
r8 37 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.135 $Y=0.157 $X2=0.135
+ $Y2=0.157
r9 36 37 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.1455 $X2=0.135 $Y2=0.157
r10 11 36 9.44419 $w=1.8e-08 $l=4.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.105 $X2=0.135 $Y2=0.1455
r11 9 35 4.64701 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.058 $X2=0.162 $Y2=0.058
r12 9 11 9.31081 $w=1.8e-08 $l=4.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.058 $X2=0.135 $Y2=0.105
r13 33 34 8.45313 $w=1.8e-08 $l=3.62e-08 $layer=M2 $thickness=3.6e-08 $X=0.216
+ $Y=0.058 $X2=0.2522 $Y2=0.058
r14 33 32 4.25571 $w=1.8e-08 $l=1.83e-08 $layer=M2 $thickness=3.6e-08 $X=0.216
+ $Y=0.058 $X2=0.1977 $Y2=0.058
r15 32 35 8.33653 $w=1.8e-08 $l=3.57e-08 $layer=M2 $thickness=3.6e-08 $X=0.1977
+ $Y=0.058 $X2=0.162 $Y2=0.058
r16 31 34 10.4352 $w=1.8e-08 $l=4.48e-08 $layer=M2 $thickness=3.6e-08 $X=0.297
+ $Y=0.058 $X2=0.2522 $Y2=0.058
r17 30 31 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.058 $X2=0.297 $Y2=0.058
r18 29 30 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.058 $X2=0.324 $Y2=0.058
r19 12 29 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.378
+ $Y=0.058 $X2=0.351 $Y2=0.058
r20 10 26 9.31081 $w=1.8e-08 $l=4.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.058 $X2=0.405 $Y2=0.105
r21 10 12 4.64701 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.058 $X2=0.378 $Y2=0.058
r22 13 26 9.44419 $w=1.8e-08 $l=4.05e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.1455 $X2=0.405 $Y2=0.105
r23 13 27 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.1455 $X2=0.405 $Y2=0.157
r24 24 27 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.405 $Y=0.157 $X2=0.405
+ $Y2=0.157
r25 8 24 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.1455 $X2=0.405 $Y2=0.157
r26 2 18 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08
+ $X=0.405 $Y=0.157 $X2=0.405 $Y2=0.157
r27 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.405
+ $Y=0.157 $X2=0.405 $Y2=0.157
r28 20 19 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.405 $Y=0.2245 $X2=0.405 $Y2=0.1755
r29 18 19 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.405 $Y=0.157 $X2=0.405 $Y2=0.1755
r30 17 18 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.405 $Y=0.1385 $X2=0.405 $Y2=0.157
r31 16 17 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.405 $Y=0.0895 $X2=0.405 $Y2=0.1385
r32 16 6 14.6259 $w=2e-08 $l=4.3e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.405 $Y=0.0895 $X2=0.405 $Y2=0.0465
.ends

.subckt PM_XOR%NET24 VSS! 6 7 3 1
c1 1 VSS! 0.00521511f $X=0.324 $Y=0.0895
c2 3 VSS! 0.00325637f $X=0.3095 $Y=0.0895
r1 7 5 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.3413 $Y=0.0895 $X2=0.3385 $Y2=0.0895
r2 1 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.324 $Y=0.0895 $X2=0.3385 $Y2=0.0895
r3 3 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.3095 $Y=0.0895 $X2=0.324 $Y2=0.0895
r4 6 3 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.3066 $Y=0.0895 $X2=0.3095 $Y2=0.0895
.ends

.subckt PM_XOR%NET27 VSS! 21 25 47 49 17 18 14 13 16 11 1 15 4 3 12 9 10
c1 1 VSS! 0.00189518f $X=0.351 $Y=0.157
c2 3 VSS! 0.00994185f $X=0.162 $Y=0.0895
c3 4 VSS! 0.0096021f $X=0.162 $Y=0.2245
c4 9 VSS! 0.042422f $X=0.351 $Y=0.0465
c5 10 VSS! 0.04493f $X=0.1475 $Y=0.0895
c6 11 VSS! 0.0450724f $X=0.1475 $Y=0.2245
c7 12 VSS! 0.0056161f $X=0.189 $Y=0.058
c8 13 VSS! 0.00545968f $X=0.189 $Y=0.256
c9 14 VSS! 0.00340201f $X=0.189 $Y=0.1845
c10 15 VSS! 0.000361978f $X=0.351 $Y=0.1455
c11 16 VSS! 0.000119895f $X=0.351 $Y=0.207
c12 17 VSS! 0.00203156f $X=0.324 $Y=0.207
c13 18 VSS! 0.000716743f $X=0.351 $Y=0.157
r1 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.1475 $Y=0.2245 $X2=0.162 $Y2=0.2245
r2 49 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.1446 $Y=0.2245 $X2=0.1475 $Y2=0.2245
r3 10 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.1475 $Y=0.0895 $X2=0.162 $Y2=0.0895
r4 47 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.1446 $Y=0.0895 $X2=0.1475 $Y2=0.0895
r5 4 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.162
+ $Y=0.2245 $X2=0.162 $Y2=0.256
r6 3 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.162
+ $Y=0.0895 $X2=0.162 $Y2=0.058
r7 44 45 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.256 $X2=0.1755 $Y2=0.256
r8 13 41 4.06646 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.256 $X2=0.189 $Y2=0.2335
r9 13 45 1.96775 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.256 $X2=0.1755 $Y2=0.256
r10 42 43 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.058 $X2=0.1755 $Y2=0.058
r11 12 38 9.77961 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.058 $X2=0.189 $Y2=0.105
r12 12 43 1.96775 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.058 $X2=0.1755 $Y2=0.058
r13 40 41 3.61444 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.218 $X2=0.189 $Y2=0.2335
r14 39 40 2.09871 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.209 $X2=0.189 $Y2=0.218
r15 37 38 12.1259 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.157 $X2=0.189 $Y2=0.105
r16 36 39 2.09871 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.209
r17 14 36 3.61444 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1845 $X2=0.189 $Y2=0.2
r18 14 37 6.41272 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1845 $X2=0.189 $Y2=0.157
r19 34 35 12.5922 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.243 $Y2=0.207
r20 34 39 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.189 $Y=0.207 $X2=0.189
+ $Y2=0.209
r21 33 35 12.5922 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.297
+ $Y=0.207 $X2=0.243 $Y2=0.207
r22 17 33 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.207 $X2=0.297 $Y2=0.207
r23 16 32 3.59766 $w=1.8e-08 $l=2.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.207 $X2=0.351 $Y2=0.1845
r24 16 17 4.64701 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.207 $X2=0.324 $Y2=0.207
r25 31 32 3.73104 $w=1.8e-08 $l=1.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.1685 $X2=0.351 $Y2=0.1845
r26 18 31 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.157 $X2=0.351 $Y2=0.1685
r27 18 29 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.351 $Y=0.157 $X2=0.351
+ $Y2=0.157
r28 15 29 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1455 $X2=0.351 $Y2=0.157
r29 1 23 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08
+ $X=0.351 $Y=0.157 $X2=0.351 $Y2=0.157
r30 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.351
+ $Y=0.157 $X2=0.351 $Y2=0.157
r31 25 24 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.351 $Y=0.2245 $X2=0.351 $Y2=0.1755
r32 23 24 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.351 $Y=0.157 $X2=0.351 $Y2=0.1755
r33 22 23 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.351 $Y=0.1385 $X2=0.351 $Y2=0.157
r34 21 22 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.351 $Y=0.0895 $X2=0.351 $Y2=0.1385
r35 21 9 14.6259 $w=2e-08 $l=4.3e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.351 $Y=0.0895 $X2=0.351 $Y2=0.0465
.ends

.subckt PM_XOR%OUT VSS! 33 19 37 48 49 11 16 17 3 15 12 1 2 10 14
c1 1 VSS! 0.00663162f $X=0.27 $Y=0.0895
c2 2 VSS! 0.00281386f $X=0.324 $Y=0.2245
c3 3 VSS! 0.00616777f $X=0.486 $Y=0.0895
c4 10 VSS! 0.0374658f $X=0.272 $Y=0.0895
c5 11 VSS! 0.0376725f $X=0.4715 $Y=0.0895
c6 12 VSS! 0.00225071f $X=0.3095 $Y=0.2245
c7 13 VSS! 0.00288649f $X=0.5135 $Y=0.058
c8 14 VSS! 0.000896201f $X=0.5135 $Y=0.211
c9 15 VSS! 0.0212155f $X=0.4725 $Y=0.058
c10 16 VSS! 0.00234455f $X=0.4995 $Y=0.211
c11 17 VSS! 0.00300856f $X=0.5135 $Y=0.105
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3413 $Y=0.2245 $X2=0.3385 $Y2=0.2245
r2 2 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.324 $Y=0.2245 $X2=0.3385 $Y2=0.2245
r3 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3095 $Y=0.2245 $X2=0.324 $Y2=0.2245
r4 48 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3066 $Y=0.2245 $X2=0.3095 $Y2=0.2245
r5 2 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.324
+ $Y=0.2245 $X2=0.324 $Y2=0.211
r6 44 45 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.211 $X2=0.3375 $Y2=0.211
r7 43 45 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.211 $X2=0.3375 $Y2=0.211
r8 42 43 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.211 $X2=0.351 $Y2=0.211
r9 41 42 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.211 $X2=0.378 $Y2=0.211
r10 40 41 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.211 $X2=0.405 $Y2=0.211
r11 39 40 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.211 $X2=0.432 $Y2=0.211
r12 38 39 5.24677 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4815
+ $Y=0.211 $X2=0.459 $Y2=0.211
r13 16 38 4.19742 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.211 $X2=0.4815 $Y2=0.211
r14 14 35 3.53581 $w=1.9e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.211 $X2=0.5135 $Y2=0.1865
r15 14 16 1.49343 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.211 $X2=0.4995 $Y2=0.211
r16 37 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.2873 $Y=0.0895 $X2=0.2845 $Y2=0.0895
r17 10 36 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.272 $Y=0.0895 $X2=0.2845 $Y2=0.0895
r18 34 35 3.83973 $w=1.9e-08 $l=1.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.1672 $X2=0.5135 $Y2=0.1865
r19 33 34 0.847733 $w=1.9e-08 $l=4.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.517
+ $Y=0.163 $X2=0.5135 $Y2=0.1672
r20 33 32 2.04453 $w=1.9e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.517
+ $Y=0.163 $X2=0.5135 $Y2=0.1527
r21 17 32 9.52453 $w=1.9e-08 $l=4.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.105 $X2=0.5135 $Y2=0.1527
r22 1 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.27
+ $Y=0.0895 $X2=0.27 $Y2=0.058
r23 13 21 1.49343 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.058 $X2=0.4995 $Y2=0.058
r24 13 17 8.02381 $w=1.9e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5135
+ $Y=0.058 $X2=0.5135 $Y2=0.105
r25 30 31 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.058 $X2=0.2835 $Y2=0.058
r26 29 31 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.058 $X2=0.2835 $Y2=0.058
r27 28 29 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.058 $X2=0.297 $Y2=0.058
r28 27 28 4.19742 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3285
+ $Y=0.058 $X2=0.3105 $Y2=0.058
r29 26 27 5.24677 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.058 $X2=0.3285 $Y2=0.058
r30 25 26 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.058 $X2=0.351 $Y2=0.058
r31 24 25 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.058 $X2=0.378 $Y2=0.058
r32 23 24 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.058 $X2=0.405 $Y2=0.058
r33 22 23 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.058 $X2=0.432 $Y2=0.058
r34 20 21 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.058 $X2=0.4995 $Y2=0.058
r35 15 20 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.058 $X2=0.486 $Y2=0.058
r36 15 22 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.058 $X2=0.459 $Y2=0.058
r37 3 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.486
+ $Y=0.0895 $X2=0.486 $Y2=0.058
r38 11 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.4715 $Y=0.0895 $X2=0.486 $Y2=0.0895
r39 19 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.4686 $Y=0.0895 $X2=0.4715 $Y2=0.0895
r40 1 10 1e-05 $l=2e-09 $X=0.27 $Y=0.0895 $X2=0.272 $Y2=0.0895
.ends

.subckt PM_XOR%A VSS! 35 16 20 49 52 12 2 1 8 7 11 13 6 5 9
c1 1 VSS! 0.00408529f $X=0.081 $Y=0.157
c2 2 VSS! 0.00222749f $X=0.459 $Y=0.157
c3 5 VSS! 0.0833987f $X=0.081 $Y=0.0465
c4 6 VSS! 0.0455271f $X=0.459 $Y=0.157
c5 7 VSS! 0.000740939f $X=0.081 $Y=0.1455
c6 8 VSS! 0.000386245f $X=0.459 $Y=0.1455
c7 9 VSS! 0.00271992f $X=0.081 $Y=0.256
c8 10 VSS! 0.00299627f $X=0.459 $Y=0.256
c9 11 VSS! 0.0036551f $X=0.081 $Y=0.1455
c10 12 VSS! 0.0236402f $X=0.108 $Y=0.256
c11 13 VSS! 0.00712929f $X=0.459 $Y=0.2315
r1 52 51 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.459 $Y=0.2245 $X2=0.459 $Y2=0.1755
r2 49 50 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.459 $Y=0.0895 $X2=0.459 $Y2=0.1385
r3 6 50 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.459 $Y=0.157 $X2=0.459 $Y2=0.1385
r4 6 51 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.459 $Y=0.157 $X2=0.459 $Y2=0.1755
r5 2 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.459
+ $Y=0.157 $X2=0.459 $Y2=0.157
r6 2 6 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08 $X=0.459
+ $Y=0.157 $X2=0.459 $Y2=0.157
r7 8 44 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1455 $X2=0.459 $Y2=0.157
r8 42 43 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.157 $X2=0.459 $Y2=0.1685
r9 42 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.459 $Y=0.157 $X2=0.459
+ $Y2=0.157
r10 40 43 5.82974 $w=1.8e-08 $l=2.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.1935 $X2=0.459 $Y2=0.1685
r11 13 40 8.86121 $w=1.8e-08 $l=3.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.2315 $X2=0.459 $Y2=0.1935
r12 10 39 4.64701 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.256 $X2=0.432 $Y2=0.256
r13 10 13 4.06404 $w=1.8e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.256 $X2=0.459 $Y2=0.2315
r14 38 39 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.256 $X2=0.432 $Y2=0.256
r15 37 38 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.378
+ $Y=0.256 $X2=0.405 $Y2=0.256
r16 36 37 21.0454 $w=1.8e-08 $l=9.03e-08 $layer=M2 $thickness=3.6e-08 $X=0.2877
+ $Y=0.256 $X2=0.378 $Y2=0.256
r17 35 36 16.9646 $w=1.8e-08 $l=7.27e-08 $layer=M2 $thickness=3.6e-08 $X=0.215
+ $Y=0.257 $X2=0.2877 $Y2=0.256
r18 35 34 4.13912 $w=1.8e-08 $l=1.78e-08 $layer=M2 $thickness=3.6e-08 $X=0.215
+ $Y=0.257 $X2=0.1972 $Y2=0.256
r19 33 34 8.21994 $w=1.8e-08 $l=3.52e-08 $layer=M2 $thickness=3.6e-08 $X=0.162
+ $Y=0.256 $X2=0.1972 $Y2=0.256
r20 32 33 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.256 $X2=0.162 $Y2=0.256
r21 12 32 6.29612 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.108
+ $Y=0.256 $X2=0.135 $Y2=0.256
r22 9 31 4.06404 $w=1.8e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.256 $X2=0.081 $Y2=0.2315
r23 9 12 4.64701 $w=1.8e-08 $l=2.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.256 $X2=0.108 $Y2=0.256
r24 30 31 5.71315 $w=1.8e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.207 $X2=0.081 $Y2=0.2315
r25 29 30 5.13017 $w=1.8e-08 $l=2.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.185 $X2=0.081 $Y2=0.207
r26 28 29 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.1715 $X2=0.081 $Y2=0.185
r27 27 28 0.699569 $w=1.8e-08 $l=3e-09 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.1685 $X2=0.081 $Y2=0.1715
r28 26 27 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.157 $X2=0.081 $Y2=0.1685
r29 11 26 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.081
+ $Y=0.1455 $X2=0.081 $Y2=0.157
r30 24 26 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.081 $Y=0.157 $X2=0.081
+ $Y2=0.157
r31 7 24 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.1455 $X2=0.081 $Y2=0.157
r32 1 18 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08
+ $X=0.081 $Y=0.157 $X2=0.081 $Y2=0.157
r33 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.081
+ $Y=0.157 $X2=0.081 $Y2=0.157
r34 20 19 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.081 $Y=0.2245 $X2=0.081 $Y2=0.1755
r35 18 19 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.081 $Y=0.157 $X2=0.081 $Y2=0.1755
r36 17 18 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.081 $Y=0.1385 $X2=0.081 $Y2=0.157
r37 16 17 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.081 $Y=0.0895 $X2=0.081 $Y2=0.1385
r38 16 5 14.6259 $w=2e-08 $l=4.3e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.081 $Y=0.0895 $X2=0.081 $Y2=0.0465
.ends

.subckt PM_XOR%NET1 VSS! 23 27 46 48 10 11 3 4 13 14 17 18 16 15 12 1 9
c1 1 VSS! 0.000487039f $X=0.297 $Y=0.157
c2 3 VSS! 0.0104954f $X=0.054 $Y=0.0895
c3 4 VSS! 0.0102216f $X=0.054 $Y=0.2245
c4 9 VSS! 0.00771738f $X=0.297 $Y=0.0465
c5 10 VSS! 0.0427025f $X=0.056 $Y=0.0895
c6 11 VSS! 0.0423204f $X=0.056 $Y=0.2245
c7 12 VSS! 0.00645871f $X=0.027 $Y=0.058
c8 13 VSS! 0.00619418f $X=0.027 $Y=0.256
c9 14 VSS! 0.0095135f $X=0.027 $Y=0.157
c10 15 VSS! 0.000245598f $X=0.297 $Y=0.1455
c11 16 VSS! 0.00318841f $X=0.027 $Y=0.1455
c12 17 VSS! 0.000676346f $X=0.297 $Y=0.1455
c13 18 VSS! 0.0128087f $X=0.027 $Y=0.157
r1 48 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.0713 $Y=0.2245 $X2=0.0685 $Y2=0.2245
r2 11 47 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.056 $Y=0.2245 $X2=0.0685 $Y2=0.2245
r3 46 45 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.0713 $Y=0.0895 $X2=0.0685 $Y2=0.0895
r4 10 45 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_48>
+ $thickness=1e-09 $X=0.056 $Y=0.0895 $X2=0.0685 $Y2=0.0895
r5 4 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.054
+ $Y=0.2245 $X2=0.054 $Y2=0.256
r6 3 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.054
+ $Y=0.0895 $X2=0.054 $Y2=0.058
r7 43 44 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.256 $X2=0.054 $Y2=0.256
r8 13 40 9.77961 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.256 $X2=0.027 $Y2=0.209
r9 13 43 1.96775 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.256 $X2=0.0405 $Y2=0.256
r10 41 42 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.058 $X2=0.054 $Y2=0.058
r11 12 39 9.77961 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.058 $X2=0.027 $Y2=0.105
r12 12 41 1.96775 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.058 $X2=0.0405 $Y2=0.058
r13 14 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.027 $Y=0.157 $X2=0.027
+ $Y2=0.157
r14 14 39 12.1259 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.157 $X2=0.027 $Y2=0.105
r15 14 40 12.1259 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.157 $X2=0.027 $Y2=0.209
r16 16 37 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.027
+ $Y=0.1455 $X2=0.027 $Y2=0.157
r17 35 36 31.4806 $w=1.8e-08 $l=1.35e-07 $layer=M3 $thickness=3.6e-08 $X=0.162
+ $Y=0.157 $X2=0.297 $Y2=0.157
r18 18 35 31.4806 $w=1.8e-08 $l=1.35e-07 $layer=M3 $thickness=3.6e-08 $X=0.027
+ $Y=0.157 $X2=0.162 $Y2=0.157
r19 18 37 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V2 $X=0.027 $Y=0.157 $X2=0.027
+ $Y2=0.157
r20 33 36 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V2 $X=0.297 $Y=0.157 $X2=0.297
+ $Y2=0.157
r21 17 33 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.297
+ $Y=0.1455 $X2=0.297 $Y2=0.157
r22 31 33 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.297 $Y=0.157 $X2=0.297
+ $Y2=0.157
r23 15 31 2.68168 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1455 $X2=0.297 $Y2=0.157
r24 1 25 6.74717 $w=2e-08 $layer=<ENCRYPTED_LAYER_23> $thickness=5.2e-08
+ $X=0.297 $Y=0.157 $X2=0.297 $Y2=0.157
r25 1 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_4> $X=0.297
+ $Y=0.157 $X2=0.297 $Y2=0.157
r26 27 26 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.297 $Y=0.2245 $X2=0.297 $Y2=0.1755
r27 25 26 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.297 $Y=0.157 $X2=0.297 $Y2=0.1755
r28 24 25 6.46262 $w=2e-08 $l=1.85e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.297 $Y=0.1385 $X2=0.297 $Y2=0.157
r29 23 24 16.6668 $w=2e-08 $l=4.9e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.297 $Y=0.0895 $X2=0.297 $Y2=0.1385
r30 23 9 14.6259 $w=2e-08 $l=4.3e-08 $layer=<ENCRYPTED_LAYER_23>
+ $thickness=5.6e-08 $X=0.297 $Y=0.0895 $X2=0.297 $Y2=0.0465
r31 4 11 1e-05 $l=2e-09 $X=0.054 $Y=0.2245 $X2=0.056 $Y2=0.2245
r32 3 10 1e-05 $l=2e-09 $X=0.054 $Y=0.0895 $X2=0.056 $Y2=0.0895
.ends

.subckt PM_XOR%NET4 VSS! 15 25 26 28 12 3 13 11 10 1 2
c1 1 VSS! 0.00673681f $X=0.27 $Y=0.2245
c2 2 VSS! 0.00684427f $X=0.378 $Y=0.2245
c3 3 VSS! 0.00940235f $X=0.486 $Y=0.2245
c4 10 VSS! 0.0369399f $X=0.272 $Y=0.2245
c5 11 VSS! 0.00336413f $X=0.3635 $Y=0.2245
c6 12 VSS! 0.0382641f $X=0.4715 $Y=0.2245
c7 13 VSS! 0.019486f $X=0.27 $Y=0.256
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.4715 $Y=0.2245 $X2=0.486 $Y2=0.2245
r2 28 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.4686 $Y=0.2245 $X2=0.4715 $Y2=0.2245
r3 26 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3953 $Y=0.2245 $X2=0.3925 $Y2=0.2245
r4 2 24 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.378 $Y=0.2245 $X2=0.3925 $Y2=0.2245
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3635 $Y=0.2245 $X2=0.378 $Y2=0.2245
r6 25 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.3606 $Y=0.2245 $X2=0.3635 $Y2=0.2245
r7 3 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.486
+ $Y=0.2245 $X2=0.486 $Y2=0.256
r8 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.378
+ $Y=0.2245 $X2=0.378 $Y2=0.256
r9 21 22 12.5922 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.256 $X2=0.486 $Y2=0.256
r10 20 21 12.5922 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.256 $X2=0.432 $Y2=0.256
r11 19 20 8.39483 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.256 $X2=0.378 $Y2=0.256
r12 18 19 7.34548 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.256 $X2=0.342 $Y2=0.256
r13 17 18 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.256 $X2=0.3105 $Y2=0.256
r14 16 17 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.256 $X2=0.297 $Y2=0.256
r15 13 16 3.14806 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.256 $X2=0.2835 $Y2=0.256
r16 1 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=<ENCRYPTED_LAYER_7> $X=0.27
+ $Y=0.2245 $X2=0.27 $Y2=0.256
r17 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.2873 $Y=0.2245 $X2=0.2845 $Y2=0.2245
r18 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=<ENCRYPTED_LAYER_49>
+ $thickness=1e-09 $X=0.272 $Y=0.2245 $X2=0.2845 $Y2=0.2245
r19 1 10 1e-05 $l=2e-09 $X=0.27 $Y=0.2245 $X2=0.272 $Y2=0.2245
.ends


* End of included file XOR.pex.netlist.pex



*
.SUBCKT XOR VSS! A VDD! B OUT
*
* VSS! VSS!
* A A
* VDD! VDD!
* B B
* OUT OUT
*
*

MM12 N_MM12_d N_MM12_g VDD! VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g VDD! VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD! VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VDD! VDD! pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM15_g VSS! VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 VSS! N_MM14_g N_MM14_s VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g N_MM8_s VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VSS! VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS! VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS! nmos_rvt L=2e-08 W=8.1e-08 nfin=3


* .include "XOR.pex.netlist.pxi"

* Start of included file XOR.pex.netlist.pxi
x_PM_XOR%NET16 VSS! N_MM4_d N_MM3_s N_NET16_3 N_NET16_1 PM_XOR%NET16
cc_1 N_NET16_3 N_A_2 0.000608874f $X=0.4175 $Y=0.0895
cc_2 N_NET16_3 N_A_6 0.0338867f $X=0.4175 $Y=0.0895
cc_3 N_NET16_3 N_B_2 0.000602083f $X=0.4175 $Y=0.0895
cc_4 N_NET16_3 N_B_6 0.0339633f $X=0.4175 $Y=0.0895
cc_5 N_NET16_1 N_OUT_15 0.000771458f $X=0.432 $Y=0.0895
cc_6 N_NET16_1 N_OUT_3 0.00475398f $X=0.432 $Y=0.0895
x_PM_XOR%B VSS! B N_MM4_g N_MM2_g N_MM14_g N_MM10_g N_B_11 N_B_2 N_B_1 N_B_8
+ N_B_7 N_B_13 N_B_6 N_B_5 N_B_12 N_B_9 N_B_10 PM_XOR%B
cc_7 N_B_11 N_A_12 0.000639405f $X=0.135 $Y=0.105
cc_8 N_B_2 N_A_2 0.00160918f $X=0.405 $Y=0.157
cc_9 N_B_1 N_A_1 0.00171664f $X=0.135 $Y=0.157
cc_10 N_B_8 N_A_8 0.00222568f $X=0.405 $Y=0.1455
cc_11 N_B_7 N_A_7 0.00244516f $X=0.135 $Y=0.1455
cc_12 N_B_11 N_A_11 0.00263834f $X=0.135 $Y=0.105
cc_13 N_B_13 N_A_13 0.00304127f $X=0.405 $Y=0.1455
cc_14 N_B_6 N_A_6 0.00330542f $X=0.405 $Y=0.0465
cc_15 N_B_5 N_A_5 0.00379483f $X=0.135 $Y=0.157
x_PM_XOR%NET24 VSS! N_MM8_s N_MM9_d N_NET24_3 N_NET24_1 PM_XOR%NET24
cc_16 N_NET24_3 N_NET1_1 0.000599484f $X=0.3095 $Y=0.0895
cc_17 N_NET24_3 N_NET1_9 0.0338642f $X=0.3095 $Y=0.0895
cc_18 N_NET24_3 N_NET27_1 0.000600955f $X=0.3095 $Y=0.0895
cc_19 N_NET24_3 N_NET27_9 0.0337954f $X=0.3095 $Y=0.0895
cc_20 N_NET24_1 N_OUT_15 0.000783679f $X=0.324 $Y=0.0895
cc_21 N_NET24_1 N_OUT_1 0.00479118f $X=0.324 $Y=0.0895
x_PM_XOR%NET27 VSS! N_MM9_g N_MM5_g N_MM14_s N_MM10_d N_NET27_17 N_NET27_18
+ N_NET27_14 N_NET27_13 N_NET27_16 N_NET27_11 N_NET27_1 N_NET27_15 N_NET27_4
+ N_NET27_3 N_NET27_12 N_NET27_9 N_NET27_10 PM_XOR%NET27
cc_22 N_NET27_17 N_A_7 0.000136945f $X=0.324 $Y=0.207
cc_23 N_NET27_18 N_A_13 0.000194361f $X=0.351 $Y=0.157
cc_24 N_NET27_17 N_A_11 0.000249643f $X=0.324 $Y=0.207
cc_25 N_NET27_18 N_A_12 0.000346497f $X=0.351 $Y=0.157
cc_26 N_NET27_14 N_A_12 0.000393547f $X=0.189 $Y=0.1845
cc_27 N_NET27_14 N_A_7 0.000568905f $X=0.189 $Y=0.1845
cc_28 N_NET27_13 N_A_12 0.000740911f $X=0.189 $Y=0.256
cc_29 N_NET27_16 N_A_12 0.000954277f $X=0.351 $Y=0.207
cc_30 N_NET27_17 N_A_12 0.0106392f $X=0.324 $Y=0.207
cc_31 N_NET27_11 N_B_5 0.0159318f $X=0.1475 $Y=0.2245
cc_32 N_NET27_14 N_B_7 0.00433437f $X=0.189 $Y=0.1845
cc_33 N_NET27_17 N_B_11 0.000624117f $X=0.324 $Y=0.207
cc_34 N_NET27_1 N_B_2 0.00164187f $X=0.351 $Y=0.157
cc_35 N_NET27_15 N_B_8 0.00225193f $X=0.351 $Y=0.1455
cc_36 N_NET27_4 N_B_5 0.001015f $X=0.162 $Y=0.2245
cc_37 N_NET27_3 N_B_1 0.0010371f $X=0.162 $Y=0.0895
cc_38 N_NET27_3 N_B_5 0.00106108f $X=0.162 $Y=0.0895
cc_39 N_NET27_14 N_B_11 0.00112639f $X=0.189 $Y=0.1845
cc_40 N_NET27_11 N_B_1 0.00150391f $X=0.1475 $Y=0.2245
cc_41 N_NET27_18 N_B_13 0.00235649f $X=0.351 $Y=0.157
cc_42 N_NET27_12 N_B_12 0.00247288f $X=0.189 $Y=0.058
cc_43 N_NET27_9 N_B_6 0.00330277f $X=0.351 $Y=0.0465
cc_44 N_NET27_10 N_B_5 0.0543598f $X=0.1475 $Y=0.0895
cc_45 N_NET27_15 N_NET1_15 0.00203584f $X=0.351 $Y=0.1455
cc_46 N_NET27_14 N_NET1_15 0.000686397f $X=0.189 $Y=0.1845
cc_47 N_NET27_17 N_NET1_15 0.000852613f $X=0.324 $Y=0.207
cc_48 N_NET27_1 N_NET1_1 0.00185055f $X=0.351 $Y=0.157
cc_49 N_NET27_18 N_NET1_17 0.00094923f $X=0.351 $Y=0.157
cc_50 N_NET27_17 N_NET1_18 0.0017186f $X=0.324 $Y=0.207
cc_51 N_NET27_9 N_NET1_9 0.00334505f $X=0.351 $Y=0.0465
cc_52 N_NET27_17 N_NET1_17 0.0061283f $X=0.324 $Y=0.207
x_PM_XOR%OUT VSS! OUT N_MM3_d N_MM8_d N_MM0_d N_MM5_d N_OUT_11 N_OUT_16 N_OUT_17
+ N_OUT_3 N_OUT_15 N_OUT_12 N_OUT_1 N_OUT_2 N_OUT_10 N_OUT_14 PM_XOR%OUT
cc_53 N_OUT_11 N_A_8 0.00036997f $X=0.4715 $Y=0.0895
cc_54 N_OUT_16 N_A_12 0.000617844f $X=0.4995 $Y=0.211
cc_55 N_OUT_17 N_A_8 0.00404674f $X=0.5135 $Y=0.105
cc_56 N_OUT_11 N_A_2 0.000896757f $X=0.4715 $Y=0.0895
cc_57 N_OUT_3 N_A_2 0.00092806f $X=0.486 $Y=0.0895
cc_58 N_OUT_3 N_A_6 0.00100888f $X=0.486 $Y=0.0895
cc_59 N_OUT_16 N_A_13 0.0014461f $X=0.4995 $Y=0.211
cc_60 N_OUT_16 N_A_8 0.00238075f $X=0.4995 $Y=0.211
cc_61 N_OUT_11 N_A_6 0.0344039f $X=0.4715 $Y=0.0895
cc_62 N_OUT_15 N_B_8 0.000314085f $X=0.4725 $Y=0.058
cc_63 N_OUT_15 N_B_10 0.000371684f $X=0.4725 $Y=0.058
cc_64 N_OUT_16 N_B_2 0.000413069f $X=0.4995 $Y=0.211
cc_65 N_OUT_15 N_B_13 0.00093422f $X=0.4725 $Y=0.058
cc_66 N_OUT_16 N_B_8 0.0021328f $X=0.4995 $Y=0.211
cc_67 N_OUT_15 N_B_12 0.00547303f $X=0.4725 $Y=0.058
cc_68 N_OUT_15 N_NET1_15 0.000439341f $X=0.4725 $Y=0.058
cc_69 N_OUT_12 N_NET1_9 0.0154454f $X=0.3095 $Y=0.2245
cc_70 N_OUT_1 N_NET1_1 0.000799389f $X=0.27 $Y=0.0895
cc_71 N_OUT_2 N_NET1_9 0.000829617f $X=0.324 $Y=0.2245
cc_72 N_OUT_1 N_NET1_9 0.00110244f $X=0.27 $Y=0.0895
cc_73 N_OUT_16 N_NET1_15 0.00119134f $X=0.4995 $Y=0.211
cc_74 N_OUT_12 N_NET1_1 0.00138651f $X=0.3095 $Y=0.2245
cc_75 N_OUT_10 N_NET1_9 0.053531f $X=0.272 $Y=0.0895
cc_76 N_OUT_12 N_NET27_16 0.00023711f $X=0.3095 $Y=0.2245
cc_77 N_OUT_16 N_NET27_15 0.00297774f $X=0.4995 $Y=0.211
cc_78 N_OUT_16 N_NET27_18 0.000296796f $X=0.4995 $Y=0.211
cc_79 N_OUT_16 N_NET27_17 0.000468769f $X=0.4995 $Y=0.211
cc_80 N_OUT_2 N_NET27_1 0.000595944f $X=0.324 $Y=0.2245
cc_81 N_OUT_1 N_NET27_9 0.000643003f $X=0.27 $Y=0.0895
cc_82 N_OUT_15 N_NET27_15 0.000675819f $X=0.4725 $Y=0.058
cc_83 N_OUT_1 N_NET27_14 0.000693638f $X=0.27 $Y=0.0895
cc_84 N_OUT_12 N_NET27_1 0.000712354f $X=0.3095 $Y=0.2245
cc_85 N_OUT_2 N_NET27_9 0.000840554f $X=0.324 $Y=0.2245
cc_86 N_OUT_12 N_NET27_9 0.0351459f $X=0.3095 $Y=0.2245
cc_87 N_OUT_17 N_NET4_13 0.000552223f $X=0.5135 $Y=0.105
cc_88 N_OUT_14 N_NET4_13 0.000575219f $X=0.5135 $Y=0.211
cc_89 N_OUT_12 N_NET4_11 0.000581385f $X=0.3095 $Y=0.2245
cc_90 N_OUT_12 N_NET4_10 0.00179117f $X=0.3095 $Y=0.2245
cc_91 N_OUT_2 N_NET4_13 0.000890118f $X=0.324 $Y=0.2245
cc_92 N_OUT_16 N_NET4_3 0.00128765f $X=0.4995 $Y=0.211
cc_93 N_OUT_2 N_NET4_2 0.00192054f $X=0.324 $Y=0.2245
cc_94 N_OUT_2 N_NET4_1 0.00446947f $X=0.324 $Y=0.2245
cc_95 N_OUT_16 N_NET4_13 0.0128405f $X=0.4995 $Y=0.211
x_PM_XOR%A VSS! A N_MM15_g N_MM12_g N_MM3_g N_MM1_g N_A_12 N_A_2 N_A_1 N_A_8
+ N_A_7 N_A_11 N_A_13 N_A_6 N_A_5 N_A_9 PM_XOR%A
x_PM_XOR%NET1 VSS! N_MM8_g N_MM0_g N_MM15_d N_MM12_d N_NET1_10 N_NET1_11
+ N_NET1_3 N_NET1_4 N_NET1_13 N_NET1_14 N_NET1_17 N_NET1_18 N_NET1_16 N_NET1_15
+ N_NET1_12 N_NET1_1 N_NET1_9 PM_XOR%NET1
cc_96 N_NET1_10 N_A_11 0.000332135f $X=0.056 $Y=0.0895
cc_97 N_NET1_11 N_A_5 0.01562f $X=0.056 $Y=0.2245
cc_98 N_NET1_3 N_A_5 0.00102514f $X=0.054 $Y=0.0895
cc_99 N_NET1_3 N_A_1 0.00104251f $X=0.054 $Y=0.0895
cc_100 N_NET1_4 N_A_5 0.00106523f $X=0.054 $Y=0.2245
cc_101 N_NET1_13 N_A_9 0.00108967f $X=0.027 $Y=0.256
cc_102 N_NET1_14 N_A_7 0.00448225f $X=0.027 $Y=0.157
cc_103 N_NET1_17 N_A_12 0.00145532f $X=0.297 $Y=0.1455
cc_104 N_NET1_11 N_A_1 0.00156322f $X=0.056 $Y=0.2245
cc_105 N_NET1_18 N_A_11 0.00238849f $X=0.027 $Y=0.157
cc_106 N_NET1_16 N_A_11 0.00383085f $X=0.027 $Y=0.1455
cc_107 N_NET1_10 N_A_5 0.0542777f $X=0.056 $Y=0.0895
cc_108 N_NET1_16 N_B_11 0.000100524f $X=0.027 $Y=0.1455
cc_109 N_NET1_18 N_B_7 0.000121909f $X=0.027 $Y=0.157
cc_110 N_NET1_15 N_B_12 0.000154321f $X=0.297 $Y=0.1455
cc_111 N_NET1_15 N_B_8 0.000173494f $X=0.297 $Y=0.1455
cc_112 N_NET1_3 N_B_7 0.000185015f $X=0.054 $Y=0.0895
cc_113 N_NET1_17 N_B_12 0.00248112f $X=0.297 $Y=0.1455
cc_114 N_NET1_14 N_B_7 0.000273693f $X=0.027 $Y=0.157
cc_115 N_NET1_17 N_B_13 0.000314175f $X=0.297 $Y=0.1455
cc_116 N_NET1_12 N_B_9 0.000589848f $X=0.027 $Y=0.058
cc_117 N_NET1_18 N_B_11 0.00539267f $X=0.027 $Y=0.157
x_PM_XOR%NET4 VSS! N_MM0_s N_MM5_s N_MM2_d N_MM1_d N_NET4_12 N_NET4_3 N_NET4_13
+ N_NET4_11 N_NET4_10 N_NET4_1 N_NET4_2 PM_XOR%NET4
cc_118 N_NET4_12 N_A_13 0.000309013f $X=0.4715 $Y=0.2245
cc_119 N_NET4_12 N_A_2 0.000689029f $X=0.4715 $Y=0.2245
cc_120 N_NET4_3 N_A_6 0.000941101f $X=0.486 $Y=0.2245
cc_121 N_NET4_13 N_A_12 0.00424546f $X=0.27 $Y=0.256
cc_122 N_NET4_12 N_A_6 0.0343897f $X=0.4715 $Y=0.2245
cc_123 N_NET4_11 N_B_2 0.000630009f $X=0.3635 $Y=0.2245
cc_124 N_NET4_11 N_B_6 0.0350023f $X=0.3635 $Y=0.2245
cc_125 N_NET4_10 N_NET1_1 0.00104406f $X=0.272 $Y=0.2245
cc_126 N_NET4_1 N_NET1_9 0.00103928f $X=0.27 $Y=0.2245
cc_127 N_NET4_10 N_NET1_9 0.0341686f $X=0.272 $Y=0.2245
cc_128 N_NET4_11 N_NET27_1 0.000861044f $X=0.3635 $Y=0.2245
cc_129 N_NET4_11 N_NET27_17 0.000434187f $X=0.3635 $Y=0.2245
cc_130 N_NET4_11 N_NET27_14 0.000551952f $X=0.3635 $Y=0.2245
cc_131 N_NET4_1 N_NET27_9 0.000623005f $X=0.27 $Y=0.2245
cc_132 N_NET4_13 N_NET27_16 0.000755959f $X=0.27 $Y=0.256
cc_133 N_NET4_2 N_NET27_9 0.000802217f $X=0.378 $Y=0.2245
cc_134 N_NET4_11 N_NET27_9 0.0347164f $X=0.3635 $Y=0.2245


* End of included file XOR.pex.netlist.pxi
.ENDS
*
